`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Student
// Engineer: Mohammad Mohsin Ahmed
// 
// Create Date: 19.02.2021 20:07:34
// Design Name: FPU
// Module Name: FPU_tb
// Project Name: Floating Point ALU
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module FPU_tb();

    reg [31:0] A,B;
    reg [1:0] operation;
    wire [31:0] ALU_output;
    wire overflow, underflow;
    FPU DUT (ALU_output ,overflow ,underflow ,A ,B ,operation);
    
    initial begin
        operation = 2'd0;   //Addition
        A = 32'b00111111100000000000000000000000;   //A=1
        B = 32'b00111111100000000000000000000000;   //B=1
        #10 B = 32'b00111111110000000000000000000000;   //B=1.5
        #10 A = 32'b10111111101000000000000000000000;   //A=-1.25
        #10 A = 32'b01000010111111100001000000000000;   //A = 127.03125
            B = 32'b01000001100001111000000000000000;   //B=16.9375
        
        operation = 2'd1;   //Subtraction
        A = 32'b00111111100000000000000000000000;   //A=1
        B = 32'b00111111100000000000000000000000;   //B=1
        #10 B = 32'b00111111110000000000000000000000;   //B=1.5
        #10 A = 32'b10111111101000000000000000000000;   //A=-1.25
        #10 A = 32'b01000010111111100001000000000000;   //A = 127.03125
            B = 32'b01000001100001111000000000000000;   //B=16.9375
        
        operation = 2'd2;   //Multiplication
        A = 32'b00111111100000000000000000000000;   //A=1
        B = 32'b00111111100000000000000000000000;   //B=1
        #10 B = 32'b00111111110000000000000000000000;   //B=1.5
        #10 A = 32'b10111111101000000000000000000000;   //A=-1.25
        #10 A = 32'b01000010111111100001000000000000;   //A = 127.03125
            B = 32'b01000001100001111000000000000000;   //B=16.9375
        
        operation = 2'd3;   //Division
        A = 32'b00111111100000000000000000000000;   //A=1
        B = 32'b00111111100000000000000000000000;   //B=1
        #10 B = 32'b00111111110000000000000000000000;   //B=1.5
        #10 A = 32'b10111111101000000000000000000000;   //A=-1.25
        #10 A = 32'b01000010111111100001000000000000;   //A = 127.03125
            B = 32'b01000001100001111000000000000000;   //B=16.9375
        
        #10 $finish;
    end    

endmodule
